module draw_string #(
    parameter string STR = "SCORE:",
    parameter START_X = 744,
    parameter START_Y = 100,
    parameter STRING_COLOR = 24'h00_00_00
  )(
    input   logic                         clk,
    input   logic [10:0]                  x, y,
    output  logic                         enable,
    output  logic [23:0]                  color
  );

  localparam END_X = START_X + STR.len()*16;
  localparam END_Y = START_Y + 32;

  assign color = STRING_COLOR;

  localparam logic [0:255][0:31][0:15] str_rom =
             {
               /*
                * code=0, hex=0x00, ascii="^@"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=1, hex=0x01, ascii="^A"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h70_0E,  /* 0111000000001110 */
               16'hE0_07,  /* 1110000000000111 */
               16'hCC_33,  /* 1100110000110011 */
               16'hCC_33,  /* 1100110000110011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hCC_33,  /* 1100110000110011 */
               16'hCE_73,  /* 1100111001110011 */
               16'hC7_E3,  /* 1100011111100011 */
               16'hC3_C3,  /* 1100001111000011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hC0_03,  /* 1100000000000011 */
               16'hE0_07,  /* 1110000000000111 */
               16'h70_0E,  /* 0111000000001110 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=2, hex=0x02, ascii="^B"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h7F_FE,  /* 0111111111111110 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF1_8F,  /* 1111000110001111 */
               16'hF8_1F,  /* 1111100000011111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h7F_FE,  /* 0111111111111110 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=3, hex=0x03, ascii="^C"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h38_70,  /* 0011100001110000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=4, hex=0x04, ascii="^D"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=5, hex=0x05, ascii="^E"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=6, hex=0x06, ascii="^F"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h7F_FE,  /* 0111111111111110 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h7F_FE,  /* 0111111111111110 */
               16'h3B_DC,  /* 0011101111011100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=7, hex=0x07, ascii="^G"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=8, hex=0x08, ascii="^H"
                */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hF8_1F,  /* 1111100000011111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hF8_1F,  /* 1111100000011111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */

               /*
                * code=9, hex=0x09, ascii="^I"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h38_1C,  /* 0011100000011100 */
               16'h30_0C,  /* 0011000000001100 */
               16'h30_0C,  /* 0011000000001100 */
               16'h30_0C,  /* 0011000000001100 */
               16'h30_0C,  /* 0011000000001100 */
               16'h38_1C,  /* 0011100000011100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=10, hex=0x0A, ascii="^J"
                */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hF8_1F,  /* 1111100000011111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hE3_C7,  /* 1110001111000111 */
               16'hC7_E3,  /* 1100011111100011 */
               16'hCF_F3,  /* 1100111111110011 */
               16'hCF_F3,  /* 1100111111110011 */
               16'hCF_F3,  /* 1100111111110011 */
               16'hCF_F3,  /* 1100111111110011 */
               16'hC7_E3,  /* 1100011111100011 */
               16'hE3_C7,  /* 1110001111000111 */
               16'hF0_0F,  /* 1111000000001111 */
               16'hF8_1F,  /* 1111100000011111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */

               /*
                * code=11, hex=0x0B, ascii="^K"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_FC,  /* 0000001111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h01_FC,  /* 0000000111111100 */
               16'h03_EC,  /* 0000001111101100 */
               16'h07_CC,  /* 0000011111001100 */
               16'h0F_8C,  /* 0000111110001100 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h7F_E0,  /* 0111111111100000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_E0,  /* 0111111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=12, hex=0x0C, ascii="^L"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=13, hex=0x0D, ascii="^M"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_0F,  /* 0000111100001111 */
               16'h0F_0F,  /* 0000111100001111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=14, hex=0x0E, ascii="^N"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FF,  /* 0011111111111111 */
               16'h3F_FF,  /* 0011111111111111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3F_FF,  /* 0011111111111111 */
               16'h3F_FF,  /* 0011111111111111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_0F,  /* 0011110000001111 */
               16'h3C_3F,  /* 0011110000111111 */
               16'h3C_3F,  /* 0011110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=15, hex=0x0F, ascii="^O"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hFB_DF,  /* 1111101111011111 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'hFC_3F,  /* 1111110000111111 */
               16'hFC_3F,  /* 1111110000111111 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'hFB_DF,  /* 1111101111011111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=16, hex=0x10, ascii="^P"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h80_00,  /* 1000000000000000 */
               16'hC0_00,  /* 1100000000000000 */
               16'hE0_00,  /* 1110000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hFE_00,  /* 1111111000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_80,  /* 1111111110000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_80,  /* 1111111110000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFE_00,  /* 1111111000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hE0_00,  /* 1110000000000000 */
               16'hC0_00,  /* 1100000000000000 */
               16'h80_00,  /* 1000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=17, hex=0x11, ascii="^Q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_04,  /* 0000000000000100 */
               16'h00_0C,  /* 0000000000001100 */
               16'h00_1C,  /* 0000000000011100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h01_FC,  /* 0000000111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h07_FC,  /* 0000011111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h07_FC,  /* 0000011111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h01_FC,  /* 0000000111111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_1C,  /* 0000000000011100 */
               16'h00_0C,  /* 0000000000001100 */
               16'h00_04,  /* 0000000000000100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=18, hex=0x12, ascii="^R"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=19, hex=0x13, ascii="^S"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=20, hex=0x14, ascii="^T"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FF,  /* 0011111111111111 */
               16'h7F_FF,  /* 0111111111111111 */
               16'hFB_CF,  /* 1111101111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hFB_CF,  /* 1111101111001111 */
               16'h7F_CF,  /* 0111111111001111 */
               16'h3F_CF,  /* 0011111111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=21, hex=0x15, ascii="^U"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=22, hex=0x16, ascii="^V"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=23, hex=0x17, ascii="^W"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=24, hex=0x18, ascii="^X"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=25, hex=0x19, ascii="^Y"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=26, hex=0x1A, ascii="^Z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_C0,  /* 0000000111000000 */
               16'h00_E0,  /* 0000000011100000 */
               16'h00_70,  /* 0000000001110000 */
               16'h00_38,  /* 0000000000111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_38,  /* 0000000000111000 */
               16'h00_70,  /* 0000000001110000 */
               16'h00_E0,  /* 0000000011100000 */
               16'h01_C0,  /* 0000000111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=27, hex=0x1B, ascii="^["
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0E_00,  /* 0000111000000000 */
               16'h1C_00,  /* 0001110000000000 */
               16'h38_00,  /* 0011100000000000 */
               16'h70_00,  /* 0111000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h70_00,  /* 0111000000000000 */
               16'h38_00,  /* 0011100000000000 */
               16'h1C_00,  /* 0001110000000000 */
               16'h0E_00,  /* 0000111000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=28, hex=0x1C, ascii="^\"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=29, hex=0x1D, ascii="^]"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h08_40,  /* 0000100001000000 */
               16'h18_60,  /* 0001100001100000 */
               16'h38_70,  /* 0011100001110000 */
               16'h78_78,  /* 0111100001111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h78_78,  /* 0111100001111000 */
               16'h38_70,  /* 0011100001110000 */
               16'h18_60,  /* 0001100001100000 */
               16'h08_40,  /* 0000100001000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=30, hex=0x1E, ascii="^^"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=31, hex=0x1F, ascii="^_"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=32, hex=0x20, ascii=" "
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=33, hex=0x21, ascii="!"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=34, hex=0x22, ascii="""
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h1C_38,  /* 0001110000111000 */
               16'h0C_30,  /* 0000110000110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=35, hex=0x23, ascii="#"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=36, hex=0x24, ascii="$"
                */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_1C,  /* 1111000000011100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'h7F_F0,  /* 0111111111110000 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hE0_3C,  /* 1110000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=37, hex=0x25, ascii="%"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h78_78,  /* 0111100001111000 */
               16'hFC_78,  /* 1111110001111000 */
               16'hCC_F0,  /* 1100110011110000 */
               16'hCC_F0,  /* 1100110011110000 */
               16'hFD_E0,  /* 1111110111100000 */
               16'h79_E0,  /* 0111100111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h1E_78,  /* 0001111001111000 */
               16'h1E_FC,  /* 0001111011111100 */
               16'h3C_CC,  /* 0011110011001100 */
               16'h3C_CC,  /* 0011110011001100 */
               16'h78_FC,  /* 0111100011111100 */
               16'h78_78,  /* 0111100001111000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=38, hex=0x26, ascii="&"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h1D_E0,  /* 0001110111100000 */
               16'h1F_C0,  /* 0001111111000000 */
               16'h3F_1C,  /* 0011111100011100 */
               16'h7F_BC,  /* 0111111110111100 */
               16'hFB_F8,  /* 1111101111111000 */
               16'hF1_F0,  /* 1111000111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_E0,  /* 1111000011100000 */
               16'hF0_E0,  /* 1111000011100000 */
               16'hF0_E0,  /* 1111000011100000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=39, hex=0x27, ascii="'"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=40, hex=0x28, ascii="("
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_70,  /* 0000000001110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_70,  /* 0000000001110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=41, hex=0x29, ascii=")"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0E_00,  /* 0000111000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0E_00,  /* 0000111000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=42, hex=0x2A, ascii="*"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h38_70,  /* 0011100001110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h38_70,  /* 0011100001110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=43, hex=0x2B, ascii="+"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=44, hex=0x2C, ascii=","
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=45, hex=0x2D, ascii="-"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=46, hex=0x2E, ascii="."
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=47, hex=0x2F, ascii="/"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h1E_00,  /* 0001111000000000 */
               16'h1E_00,  /* 0001111000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h78_00,  /* 0111100000000000 */
               16'h78_00,  /* 0111100000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=48, hex=0x30, ascii="0"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=49, hex=0x31, ascii="1"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_C0,  /* 0001111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=50, hex=0x32, ascii="2"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hE0_3C,  /* 1110000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=51, hex=0x33, ascii="3"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_78,  /* 0000000001111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=52, hex=0x34, ascii="4"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h07_F0,  /* 0000011111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h3E_F0,  /* 0011111011110000 */
               16'h7C_F0,  /* 0111110011110000 */
               16'hF8_F0,  /* 1111100011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h03_FC,  /* 0000001111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=53, hex=0x35, ascii="5"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=54, hex=0x36, ascii="6"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=55, hex=0x37, ascii="7"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=56, hex=0x38, ascii="8"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h78_78,  /* 0111100001111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h78_78,  /* 0111100001111000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=57, hex=0x39, ascii="9"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_FC,  /* 0111111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=58, hex=0x3A, ascii=":"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=59, hex=0x3B, ascii=";"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=60, hex=0x3C, ascii="<"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_F8,  /* 0000000011111000 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=61, hex=0x3D, ascii="="
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=62, hex=0x3E, ascii=">"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_F8,  /* 0000000011111000 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=63, hex=0x3F, ascii="?"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=64, hex=0x40, ascii="@"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF1_FC,  /* 1111000111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF1_F0,  /* 1111000111110000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'h7F_F0,  /* 0111111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=65, hex=0x41, ascii="A"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=66, hex=0x42, ascii="B"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'hFF_F8,  /* 1111111111111000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=67, hex=0x43, ascii="C"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h7C_7C,  /* 0111110001111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hF0_1C,  /* 1111000000011100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_1C,  /* 1111000000011100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'h7C_7C,  /* 0111110001111100 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=68, hex=0x44, ascii="D"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_E0,  /* 1111111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hFF_E0,  /* 1111111111100000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=69, hex=0x45, ascii="E"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_1C,  /* 0011110000011100 */
               16'h3C_0C,  /* 0011110000001100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_0C,  /* 0011110000001100 */
               16'h3C_1C,  /* 0011110000011100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=70, hex=0x46, ascii="F"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_1C,  /* 0011110000011100 */
               16'h3C_0C,  /* 0011110000001100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_C0,  /* 0011110011000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=71, hex=0x47, ascii="G"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h7C_7C,  /* 0111110001111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hF0_1C,  /* 1111000000011100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF1_FC,  /* 1111000111111100 */
               16'hF1_FC,  /* 1111000111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'h7C_7C,  /* 0111110001111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_EC,  /* 0001111111101100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=72, hex=0x48, ascii="H"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=73, hex=0x49, ascii="I"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=74, hex=0x4A, ascii="J"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_FC,  /* 0000001111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_E0,  /* 0111111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=75, hex=0x4B, ascii="K"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3D_F0,  /* 0011110111110000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3D_F0,  /* 0011110111110000 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=76, hex=0x4C, ascii="L"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_0C,  /* 0011110000001100 */
               16'h3C_1C,  /* 0011110000011100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=77, hex=0x4D, ascii="M"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hFC_FC,  /* 1111110011111100 */
               16'hFC_FC,  /* 1111110011111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=78, hex=0x4E, ascii="N"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFE_3C,  /* 1111111000111100 */
               16'hFE_3C,  /* 1111111000111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF1_FC,  /* 1111000111111100 */
               16'hF1_FC,  /* 1111000111111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_7C,  /* 1111000001111100 */
               16'hF0_7C,  /* 1111000001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=79, hex=0x4F, ascii="O"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=80, hex=0x50, ascii="P"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=81, hex=0x51, ascii="Q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_BC,  /* 1111001110111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF9_FC,  /* 1111100111111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_E0,  /* 0000000011100000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=82, hex=0x52, ascii="R"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3D_F0,  /* 0011110111110000 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=83, hex=0x53, ascii="S"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'h78_00,  /* 0111100000000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=84, hex=0x54, ascii="T"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hC7_8C,  /* 1100011110001100 */
               16'hC7_8C,  /* 1100011110001100 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=85, hex=0x55, ascii="U"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=86, hex=0x56, ascii="V"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=87, hex=0x57, ascii="W"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h38_70,  /* 0011100001110000 */
               16'h38_70,  /* 0011100001110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=88, hex=0x58, ascii="X"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h78_78,  /* 0111100001111000 */
               16'h78_78,  /* 0111100001111000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h78_78,  /* 0111100001111000 */
               16'h78_78,  /* 0111100001111000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=89, hex=0x59, ascii="Y"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=90, hex=0x5A, ascii="Z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hE0_3C,  /* 1110000000111100 */
               16'hC0_3C,  /* 1100000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_1C,  /* 1111000000011100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=91, hex=0x5B, ascii="["
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=92, hex=0x5C, ascii="\"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h78_00,  /* 0111100000000000 */
               16'h78_00,  /* 0111100000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h1E_00,  /* 0001111000000000 */
               16'h1E_00,  /* 0001111000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_78,  /* 0000000001111000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=93, hex=0x5D, ascii="]"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=94, hex=0x5E, ascii="^"
                */
               16'h03_00,  /* 0000001100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h78_78,  /* 0111100001111000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hE0_1C,  /* 1110000000011100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=95, hex=0x5F, ascii="_"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=96, hex=0x60, ascii="`"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=97, hex=0x61, ascii="a"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F0,  /* 0111111111110000 */
               16'hF8_F0,  /* 1111100011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_FC,  /* 0111111111111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=98, hex=0x62, ascii="b"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3F_80,  /* 0011111110000000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=99, hex=0x63, ascii="c"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=100, hex=0x64, ascii="d"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h1F_F0,  /* 0001111111110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h78_F0,  /* 0111100011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h79_F0,  /* 0111100111110000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h1F_3C,  /* 0001111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=101, hex=0x65, ascii="e"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=102, hex=0x66, ascii="f"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_70,  /* 0011110001110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=103, hex=0x67, ascii="g"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h7F_FC,  /* 0111111111111100 */
               16'hF9_F0,  /* 1111100111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF8_F0,  /* 1111100011110000 */
               16'h7F_F0,  /* 0111111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_E0,  /* 0111111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=104, hex=0x68, ascii="h"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=105, hex=0x69, ascii="i"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_80,  /* 0001111110000000 */
               16'h1F_80,  /* 0001111110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=106, hex=0x6A, ascii="j"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=107, hex=0x6B, ascii="k"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'hFC_00,  /* 1111110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3D_F0,  /* 0011110111110000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_E0,  /* 0011111111100000 */
               16'h3D_F0,  /* 0011110111110000 */
               16'h3C_F8,  /* 0011110011111000 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=108, hex=0x6C, ascii="l"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h1F_80,  /* 0001111110000000 */
               16'h1F_80,  /* 0001111110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=109, hex=0x6D, ascii="m"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFC_F0,  /* 1111110011110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=110, hex=0x6E, ascii="n"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=111, hex=0x6F, ascii="o"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=112, hex=0x70, ascii="p"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_7C,  /* 0011110001111100 */
               16'h3F_F8,  /* 0011111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=113, hex=0x71, ascii="q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h7F_FC,  /* 0111111111111100 */
               16'hF9_F0,  /* 1111100111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF8_F0,  /* 1111100011110000 */
               16'h7F_F0,  /* 0111111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h03_FC,  /* 0000001111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=114, hex=0x72, ascii="r"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hFF_F8,  /* 1111111111111000 */
               16'h3F_7C,  /* 0011111101111100 */
               16'h3E_3C,  /* 0011111000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=115, hex=0x73, ascii="s"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'hF0_7C,  /* 1111000001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h78_00,  /* 0111100000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_80,  /* 0001111110000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_78,  /* 0000000001111000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=116, hex=0x74, ascii="t"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_00,  /* 0000000100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h07_00,  /* 0000011100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_1C,  /* 0000111100011100 */
               16'h0F_BC,  /* 0000111110111100 */
               16'h07_F8,  /* 0000011111111000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=117, hex=0x75, ascii="u"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'h7F_FC,  /* 0111111111111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=118, hex=0x76, ascii="v"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3E_7C,  /* 0011111001111100 */
               16'h1F_F8,  /* 0001111111111000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_80,  /* 0000000110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=119, hex=0x77, ascii="w"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF3_3C,  /* 1111001100111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hF7_BC,  /* 1111011110111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h38_70,  /* 0011100001110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=120, hex=0x78, ascii="x"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7C_F8,  /* 0111110011111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=121, hex=0x79, ascii="y"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'h7F_FC,  /* 0111111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_7C,  /* 0000000001111100 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'hFF_E0,  /* 1111111111100000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=122, hex=0x7A, ascii="z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_F8,  /* 1111000011111000 */
               16'hF1_F0,  /* 1111000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=123, hex=0x7B, ascii="{"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_FC,  /* 0000000011111100 */
               16'h01_FC,  /* 0000000111111100 */
               16'h03_E0,  /* 0000001111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h01_FC,  /* 0000000111111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=124, hex=0x7C, ascii="|"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=125, hex=0x7D, ascii="}"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_80,  /* 0011111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h01_E0,  /* 0000000111100000 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h01_E0,  /* 0000000111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h3F_80,  /* 0011111110000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=126, hex=0x7E, ascii="~"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_1C,  /* 0011110000011100 */
               16'h7F_3C,  /* 0111111100111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF3_F8,  /* 1111001111111000 */
               16'hE0_F0,  /* 1110000011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=127, hex=0x7F, ascii="^?"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h7C_F8,  /* 0111110011111000 */
               16'hF8_7C,  /* 1111100001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=128, hex=0x80, ascii="!^@"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_0C,  /* 1111000000001100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=129, hex=0x81, ascii="!^A"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=130, hex=0x82, ascii="!^B"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=131, hex=0x83, ascii="!^C"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=132, hex=0x84, ascii="!^D"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=133, hex=0x85, ascii="!^E"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=134, hex=0x86, ascii="!^F"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=135, hex=0x87, ascii="!^G"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=136, hex=0x88, ascii="!^H"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=137, hex=0x89, ascii="!^I"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=138, hex=0x8A, ascii="!^J"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=139, hex=0x8B, ascii="!^K"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=140, hex=0x8C, ascii="!^L"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=141, hex=0x8D, ascii="!^M"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=142, hex=0x8E, ascii="!^N"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=143, hex=0x8F, ascii="!^O"
                */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=144, hex=0x90, ascii="!^P"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=145, hex=0x91, ascii="!^Q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'h3C_FC,  /* 0011110011111100 */
               16'h3C_FC,  /* 0011110011111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=146, hex=0x92, ascii="!^R"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=147, hex=0x93, ascii="!^S"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h03_00,  /* 0000001100000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=148, hex=0x94, ascii="!^T"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=149, hex=0x95, ascii="!^U"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=150, hex=0x96, ascii="!^V"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=151, hex=0x97, ascii="!^W"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=152, hex=0x98, ascii="!^X"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=153, hex=0x99, ascii="!^Y"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=154, hex=0x9A, ascii="!^Z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=155, hex=0x9B, ascii="!^["
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=156, hex=0x9C, ascii="!^\"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_30,  /* 0011110000110000 */
               16'h3C_30,  /* 0011110000110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFF_F0,  /* 1111111111110000 */
               16'hFF_F0,  /* 1111111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=157, hex=0x9D, ascii="!^]"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=158, hex=0x9E, ascii="!^^"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hF0_30,  /* 1111000000110000 */
               16'hF0_30,  /* 1111000000110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=159, hex=0x9F, ascii="!^_"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_FC,  /* 0000000011111100 */
               16'h00_FC,  /* 0000000011111100 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=160, hex=0xA0, ascii="! "
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=161, hex=0xA1, ascii="!!"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=162, hex=0xA2, ascii="!""
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=163, hex=0xA3, ascii="!#"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=164, hex=0xA4, ascii="!$"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=165, hex=0xA5, ascii="!%"
                */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFC_3C,  /* 1111110000111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF3_FC,  /* 1111001111111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=166, hex=0xA6, ascii="!&"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=167, hex=0xA7, ascii="!'"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=168, hex=0xA8, ascii="!("
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_00,  /* 1111100000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_7C,  /* 1111100001111100 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=169, hex=0xA9, ascii="!)"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=170, hex=0xAA, ascii="!*"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=171, hex=0xAB, ascii="!+"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hC0_3C,  /* 1100000000111100 */
               16'hC0_3C,  /* 1100000000111100 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=172, hex=0xAC, ascii="!,"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_0C,  /* 1111000000001100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hF0_FC,  /* 1111000011111100 */
               16'hC3_FC,  /* 1100001111111100 */
               16'hC3_FC,  /* 1100001111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=173, hex=0xAD, ascii="!-"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h07_E0,  /* 0000011111100000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=174, hex=0xAE, ascii="!."
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0E_1C,  /* 0000111000011100 */
               16'h1E_3C,  /* 0001111000111100 */
               16'h3C_78,  /* 0011110001111000 */
               16'h78_F0,  /* 0111100011110000 */
               16'hF1_E0,  /* 1111000111100000 */
               16'hF1_E0,  /* 1111000111100000 */
               16'h78_F0,  /* 0111100011110000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h1E_3C,  /* 0001111000111100 */
               16'h0E_1C,  /* 0000111000011100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=175, hex=0xAF, ascii="!/"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hE1_C0,  /* 1110000111000000 */
               16'hF1_E0,  /* 1111000111100000 */
               16'h78_F0,  /* 0111100011110000 */
               16'h3C_78,  /* 0011110001111000 */
               16'h1E_3C,  /* 0001111000111100 */
               16'h1E_3C,  /* 0001111000111100 */
               16'h3C_78,  /* 0011110001111000 */
               16'h78_F0,  /* 0111100011110000 */
               16'hF1_E0,  /* 1111000111100000 */
               16'hE1_C0,  /* 1110000111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=176, hex=0xB0, ascii="!0"
                */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */
               16'h03_03,  /* 0000001100000011 */
               16'h03_03,  /* 0000001100000011 */
               16'h30_30,  /* 0011000000110000 */
               16'h30_30,  /* 0011000000110000 */

               /*
                * code=177, hex=0xB1, ascii="!1"
                */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */
               16'h33_33,  /* 0011001100110011 */
               16'h33_33,  /* 0011001100110011 */
               16'hCC_CC,  /* 1100110011001100 */
               16'hCC_CC,  /* 1100110011001100 */

               /*
                * code=178, hex=0xB2, ascii="!2"
                */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */
               16'hF3_F3,  /* 1111001111110011 */
               16'hF3_F3,  /* 1111001111110011 */
               16'h3F_3F,  /* 0011111100111111 */
               16'h3F_3F,  /* 0011111100111111 */

               /*
                * code=179, hex=0xB3, ascii="!3"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=180, hex=0xB4, ascii="!4"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=181, hex=0xB5, ascii="!5"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=182, hex=0xB6, ascii="!6"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=183, hex=0xB7, ascii="!7"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=184, hex=0xB8, ascii="!8"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=185, hex=0xB9, ascii="!9"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=186, hex=0xBA, ascii="!:"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=187, hex=0xBB, ascii="!;"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=188, hex=0xBC, ascii="!<"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'hFF_3C,  /* 1111111100111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=189, hex=0xBD, ascii="!="
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=190, hex=0xBE, ascii="!>"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=191, hex=0xBF, ascii="!?"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=192, hex=0xC0, ascii="!@"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=193, hex=0xC1, ascii="!A"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=194, hex=0xC2, ascii="!B"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=195, hex=0xC3, ascii="!C"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=196, hex=0xC4, ascii="!D"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=197, hex=0xC5, ascii="!E"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=198, hex=0xC6, ascii="!F"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=199, hex=0xC7, ascii="!G"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=200, hex=0xC8, ascii="!H"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=201, hex=0xC9, ascii="!I"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=202, hex=0xCA, ascii="!J"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_3F,  /* 1111111100111111 */
               16'hFF_3F,  /* 1111111100111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=203, hex=0xCB, ascii="!K"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_3F,  /* 1111111100111111 */
               16'hFF_3F,  /* 1111111100111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=204, hex=0xCC, ascii="!L"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3F,  /* 0000111100111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=205, hex=0xCD, ascii="!M"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=206, hex=0xCE, ascii="!N"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_3F,  /* 1111111100111111 */
               16'hFF_3F,  /* 1111111100111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_3F,  /* 1111111100111111 */
               16'hFF_3F,  /* 1111111100111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=207, hex=0xCF, ascii="!O"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=208, hex=0xD0, ascii="!P"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=209, hex=0xD1, ascii="!Q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=210, hex=0xD2, ascii="!R"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=211, hex=0xD3, ascii="!S"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=212, hex=0xD4, ascii="!T"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=213, hex=0xD5, ascii="!U"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=214, hex=0xD6, ascii="!V"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_FF,  /* 0000111111111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=215, hex=0xD7, ascii="!W"
                */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */
               16'h0F_3C,  /* 0000111100111100 */

               /*
                * code=216, hex=0xD8, ascii="!X"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=217, hex=0xD9, ascii="!Y"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=218, hex=0xDA, ascii="!Z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_FF,  /* 0000001111111111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=219, hex=0xDB, ascii="!["
                */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */

               /*
                * code=220, hex=0xDC, ascii="!\"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */

               /*
                * code=221, hex=0xDD, ascii="!]"
                */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */
               16'hFF_00,  /* 1111111100000000 */

               /*
                * code=222, hex=0xDE, ascii="!^"
                */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */

               /*
                * code=223, hex=0xDF, ascii="!_"
                */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'hFF_FF,  /* 1111111111111111 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=224, hex=0xE0, ascii="!`"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=225, hex=0xE1, ascii="!a"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_C0,  /* 0011111111000000 */
               16'h7F_E0,  /* 0111111111100000 */
               16'hF9_F0,  /* 1111100111110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'hF1_E0,  /* 1111000111100000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_E0,  /* 1111001111100000 */
               16'hF1_F0,  /* 1111000111110000 */
               16'hF0_F8,  /* 1111000011111000 */
               16'hF0_7C,  /* 1111000001111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_7C,  /* 1111000001111100 */
               16'hF0_F8,  /* 1111000011111000 */
               16'hF0_F0,  /* 1111000011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=226, hex=0xE2, ascii="!b"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=227, hex=0xE3, ascii="!c"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=228, hex=0xE4, ascii="!d"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF8_3C,  /* 1111100000111100 */
               16'h7C_00,  /* 0111110000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'hF8_3C,  /* 1111100000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=229, hex=0xE5, ascii="!e"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=230, hex=0xE6, ascii="!f"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=231, hex=0xE7, ascii="!g"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=232, hex=0xE8, ascii="!h"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=233, hex=0xE9, ascii="!i"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=234, hex=0xEA, ascii="!j"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'hFC_FC,  /* 1111110011111100 */
               16'hFC_FC,  /* 1111110011111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=235, hex=0xEB, ascii="!k"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_FC,  /* 0000001111111100 */
               16'h03_FC,  /* 0000001111111100 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h0F_FC,  /* 0000111111111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h3C_3C,  /* 0011110000111100 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=236, hex=0xEC, ascii="!l"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=237, hex=0xED, ascii="!m"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_0F,  /* 0000000000001111 */
               16'h00_0F,  /* 0000000000001111 */
               16'h00_3C,  /* 0000000000111100 */
               16'h00_3C,  /* 0000000000111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hF3_CF,  /* 1111001111001111 */
               16'hFF_0F,  /* 1111111100001111 */
               16'hFF_0F,  /* 1111111100001111 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3F_FC,  /* 0011111111111100 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'hF0_00,  /* 1111000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=238, hex=0xEE, ascii="!n"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=239, hex=0xEF, ascii="!o"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'hF0_3C,  /* 1111000000111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=240, hex=0xF0, ascii="!p"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=241, hex=0xF1, ascii="!q"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=242, hex=0xF2, ascii="!r"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_F8,  /* 0000000011111000 */
               16'h00_F8,  /* 0000000011111000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=243, hex=0xF3, ascii="!s"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'h7C_00,  /* 0111110000000000 */
               16'h3E_00,  /* 0011111000000000 */
               16'h1F_00,  /* 0001111100000000 */
               16'h0F_80,  /* 0000111110000000 */
               16'h07_C0,  /* 0000011111000000 */
               16'h03_E0,  /* 0000001111100000 */
               16'h01_F0,  /* 0000000111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h7F_F8,  /* 0111111111111000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=244, hex=0xF4, ascii="!t"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_FC,  /* 0000000011111100 */
               16'h01_FE,  /* 0000000111111110 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_CF,  /* 0000001111001111 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */

               /*
                * code=245, hex=0xF5, ascii="!u"
                */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'h7F_80,  /* 0111111110000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=246, hex=0xF6, ascii="!v"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'hFF_FC,  /* 1111111111111100 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h07_80,  /* 0000011110000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=247, hex=0xF7, ascii="!w"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_3C,  /* 0011111100111100 */
               16'h3F_3C,  /* 0011111100111100 */
               16'hF3_F0,  /* 1111001111110000 */
               16'hF3_F0,  /* 1111001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=248, hex=0xF8, ascii="!x"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h1F_E0,  /* 0001111111100000 */
               16'h0F_C0,  /* 0000111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=249, hex=0xF9, ascii="!y"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=250, hex=0xFA, ascii="!z"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h03_C0,  /* 0000001111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=251, hex=0xFB, ascii="!{"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_FF,  /* 0000000011111111 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'h00_F0,  /* 0000000011110000 */
               16'hFC_F0,  /* 1111110011110000 */
               16'hFC_F0,  /* 1111110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h0F_F0,  /* 0000111111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h03_F0,  /* 0000001111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=252, hex=0xFC, ascii="!|"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF7_E0,  /* 1111011111100000 */
               16'h3E_F0,  /* 0011111011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h3C_F0,  /* 0011110011110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=253, hex=0xFD, ascii="!}"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'h3F_00,  /* 0011111100000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'hF3_C0,  /* 1111001111000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h0F_00,  /* 0000111100000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'h3C_00,  /* 0011110000000000 */
               16'hF0_C0,  /* 1111000011000000 */
               16'hF0_C0,  /* 1111000011000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'hFF_C0,  /* 1111111111000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=254, hex=0xFE, ascii="!~"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h3F_F0,  /* 0011111111110000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */

               /*
                * code=255, hex=0xFF, ascii="!^"
                */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00,  /* 0000000000000000 */
               16'h00_00   /* 0000000000000000 */
             };

  logic [0:STR.len()-1][0:31][0:15] disp;
  integer i,j;

  always_comb
    begin
      for (i = 0; i < STR.len(); ++i)
        begin
          disp [i] = str_rom[STR.getc(i)];
        end
    end

  always_ff @(posedge clk)
    begin
      if (x >= START_X && x < END_X
          && y >=START_Y && y < END_Y)
        enable <= disp[(x - START_X) / 16][(y - START_Y) % 32][(x - START_X) % 16];
      else
        enable <= 0;
    end
endmodule
