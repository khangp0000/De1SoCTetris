module draw_number #(
    parameter NUM_DISPLAY = 8,
    parameter INPUT_WIDTH = 27,
    parameter START_X = 840,
    parameter START_Y = 100,
    parameter NUM_COLOR = 24'h00_00_00
  )(
    input   logic                         clk,
    input   logic [10:0]                  x, y,
    input   logic [INPUT_WIDTH - 1 : 0]   in,
    output  logic                         enable,
    output  logic [23:0]                  color
  );

  localparam END_X = START_X + NUM_DISPLAY*16;
  localparam END_Y = START_Y + 32;

  assign color = NUM_COLOR;

  // logic [0:NUM_DISPLAY - 1][0:32][0:16] disp;
  logic [0:NUM_DISPLAY - 1][3:0] number_to_display;

  integer i,j;

  logic [0:9][0:31][0:15] rom =
        {
          /*
           * ascii="0"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h1F_E0,  /* 0001111111100000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h7C_F8,  /* 0111110011111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF3_3C,  /* 1111001100111100 */
          16'hF7_BC,  /* 1111011110111100 */
          16'hF7_BC,  /* 1111011110111100 */
          16'hF7_BC,  /* 1111011110111100 */
          16'hF7_BC,  /* 1111011110111100 */
          16'hF3_3C,  /* 1111001100111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7C_F8,  /* 0111110011111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h1F_E0,  /* 0001111111100000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="1"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h07_C0,  /* 0000011111000000 */
          16'h0F_C0,  /* 0000111111000000 */
          16'h1F_C0,  /* 0001111111000000 */
          16'h3F_C0,  /* 0011111111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h03_C0,  /* 0000001111000000 */
          16'h3F_FC,  /* 0011111111111100 */
          16'h3F_FC,  /* 0011111111111100 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="2"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h7F_F8,  /* 0111111111111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hE0_3C,  /* 1110000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_7C,  /* 0000000001111100 */
          16'h00_F8,  /* 0000000011111000 */
          16'h01_F0,  /* 0000000111110000 */
          16'h03_E0,  /* 0000001111100000 */
          16'h07_C0,  /* 0000011111000000 */
          16'h0F_80,  /* 0000111110000000 */
          16'h1F_00,  /* 0001111100000000 */
          16'h3E_00,  /* 0011111000000000 */
          16'h7C_00,  /* 0111110000000000 */
          16'hF8_00,  /* 1111100000000000 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hFF_FC,  /* 1111111111111100 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="3"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h7F_F8,  /* 0111111111111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_78,  /* 0000000001111000 */
          16'h0F_F0,  /* 0000111111110000 */
          16'h0F_F0,  /* 0000111111110000 */
          16'h00_78,  /* 0000000001111000 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7F_F8,  /* 0111111111111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="4"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h01_F0,  /* 0000000111110000 */
          16'h03_F0,  /* 0000001111110000 */
          16'h07_F0,  /* 0000011111110000 */
          16'h0F_F0,  /* 0000111111110000 */
          16'h1F_F0,  /* 0001111111110000 */
          16'h3E_F0,  /* 0011111011110000 */
          16'h7C_F0,  /* 0111110011110000 */
          16'hF8_F0,  /* 1111100011110000 */
          16'hF0_F0,  /* 1111000011110000 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hFF_FC,  /* 1111111111111100 */
          16'h00_F0,  /* 0000000011110000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h00_F0,  /* 0000000011110000 */
          16'h03_FC,  /* 0000001111111100 */
          16'h03_FC,  /* 0000001111111100 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="5"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hFF_F0,  /* 1111111111110000 */
          16'hFF_F8,  /* 1111111111111000 */
          16'h00_7C,  /* 0000000001111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7F_F8,  /* 0111111111111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="6"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h0F_F0,  /* 0000111111110000 */
          16'h1F_F0,  /* 0001111111110000 */
          16'h3E_00,  /* 0011111000000000 */
          16'h7C_00,  /* 0111110000000000 */
          16'hF8_00,  /* 1111100000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hF0_00,  /* 1111000000000000 */
          16'hFF_F0,  /* 1111111111110000 */
          16'hFF_F8,  /* 1111111111111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7F_F8,  /* 0111111111111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="7"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hFF_FC,  /* 1111111111111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_7C,  /* 0000000001111100 */
          16'h00_F8,  /* 0000000011111000 */
          16'h01_F0,  /* 0000000111110000 */
          16'h03_E0,  /* 0000001111100000 */
          16'h07_C0,  /* 0000011111000000 */
          16'h0F_80,  /* 0000111110000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h0F_00,  /* 0000111100000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="8"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h7F_F8,  /* 0111111111111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'h78_78,  /* 0111100001111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h78_78,  /* 0111100001111000 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7F_F8,  /* 0111111111111000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */

          /*
           * ascii="9"
           */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h3F_F0,  /* 0011111111110000 */
          16'h7F_F8,  /* 0111111111111000 */
          16'hF8_7C,  /* 1111100001111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF0_3C,  /* 1111000000111100 */
          16'hF8_7C,  /* 1111100001111100 */
          16'h7F_FC,  /* 0111111111111100 */
          16'h3F_FC,  /* 0011111111111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_3C,  /* 0000000000111100 */
          16'h00_7C,  /* 0000000001111100 */
          16'h00_F8,  /* 0000000011111000 */
          16'h01_F0,  /* 0000000111110000 */
          16'h3F_E0,  /* 0011111111100000 */
          16'h3F_C0,  /* 0011111111000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00,  /* 0000000000000000 */
          16'h00_00   /* 0000000000000000 */
        };

  always_comb
    begin
      for (i = 0; i < NUM_DISPLAY; ++i)
        begin
          number_to_display[NUM_DISPLAY - 1 - i] = in/(10**i)%10;
        end
    end

  // always_ff @(posedge clk) // NUM_DISPLAY port ROM ?
  //   begin
  //     for (j = 0; j < NUM_DISPLAY; ++j)
  //       begin
  //         disp[j] <<= rom[number_to_display[j]];
  //       end
  //   end

  always_ff @(posedge clk)
    begin
      if (x >= START_X && x < END_X
          && y >=START_Y && y < END_Y)
        enable <= rom[number_to_display[(x - START_X) / 16]][(y - START_Y) % 32][(x - START_X) % 16];
      else
        enable <= 0;
    end

endmodule 
